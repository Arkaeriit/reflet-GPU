/*------------------------------------\
|ROM containing the font Public Pixel.|
|Made by GGBotNet under the license   |
|Creative Commons Zero v1.0 Universal.|
|Accepts ISO/IEC 8859-1 encoded       |
|characters as input.                 |
\------------------------------------*/

module public_pixel (
    input [7:0] char,
    input [$clog2(64)-1:0] index,
    output is_foreground
    );

    reg [63:0] font_char;
    wire [63:0] shift = font_char >> index;
    assign is_foreground = shift[0];
    
    always @ (char)
        case(char)
            8'h21 : font_char = 64'h0C000C1E1E1E0C00;
            8'h22 : font_char = 64'h0000001224363600;
            8'h23 : font_char = 64'h367F3636367F3600;
            8'h24 : font_char = 64'h083F683E0B7E0800;
            8'h25 : font_char = 64'h23562C1832654200;
            8'h26 : font_char = 64'h3E63735B0E1B0E00;
            8'h27 : font_char = 64'h00000004080C0C00;
            8'h28 : font_char = 64'h380C0606060C3800;
            8'h29 : font_char = 64'h0E18303030180E00;
            8'h2A : font_char = 64'h00000000361C3600;
            8'h2B : font_char = 64'h08083E0808000000;
            8'h2C : font_char = 64'h04080C0C00000000;
            8'h2D : font_char = 64'h00003E0000000000;
            8'h2E : font_char = 64'h0C0C000000000000;
            8'h2F : font_char = 64'h0103060C18302000;
            8'h30 : font_char = 64'h3E67636363733E00;
            8'h31 : font_char = 64'h7E18181818181E00;
            8'h32 : font_char = 64'h7F03061C30633E00;
            8'h33 : font_char = 64'h3E63603C60633E00;
            8'h34 : font_char = 64'h60607F63666C7800;
            8'h35 : font_char = 64'h3E6360603F037F00;
            8'h36 : font_char = 64'h3E63633F03633E00;
            8'h37 : font_char = 64'h03060C1830637F00;
            8'h38 : font_char = 64'h3E63633E63633E00;
            8'h39 : font_char = 64'h3E63607E63633E00;
            8'h3A : font_char = 64'h0C0C000C0C000000;
            8'h3B : font_char = 64'h080C000C0C000000;
            8'h3C : font_char = 64'h381C0E1C38000000;
            8'h3D : font_char = 64'h003E003E00000000;
            8'h3E : font_char = 64'h0E1C381C0E000000;
            8'h3F : font_char = 64'h0C000C3C60633E00;
            8'h40 : font_char = 64'h3E033B6B6B633E00;
            8'h41 : font_char = 64'h63637F6363361C00;
            8'h42 : font_char = 64'h3F63633F63633F00;
            8'h43 : font_char = 64'h3E63030303633E00;
            8'h44 : font_char = 64'h1F33636363331F00;
            8'h45 : font_char = 64'h7F03031F03037F00;
            8'h46 : font_char = 64'h0303031F03037F00;
            8'h47 : font_char = 64'h7E63637B03037E00;
            8'h48 : font_char = 64'h6363637F63636300;
            8'h49 : font_char = 64'h7E18181818187E00;
            8'h4A : font_char = 64'h3E63636060607800;
            8'h4B : font_char = 64'h63331B0F1B336300;
            8'h4C : font_char = 64'h7F03030303030300;
            8'h4D : font_char = 64'h6363636B7F776300;
            8'h4E : font_char = 64'h6363737B6F676300;
            8'h4F : font_char = 64'h3E63636363633E00;
            8'h50 : font_char = 64'h0303033F63633F00;
            8'h51 : font_char = 64'h5E337B6363633E00;
            8'h52 : font_char = 64'h63331B3F63633F00;
            8'h53 : font_char = 64'h3E63603E03633E00;
            8'h54 : font_char = 64'h1818181818187E00;
            8'h55 : font_char = 64'h3E63636363636300;
            8'h56 : font_char = 64'h081C366363636300;
            8'h57 : font_char = 64'h6363777F6B636300;
            8'h58 : font_char = 64'h63773E1C3E776300;
            8'h59 : font_char = 64'h1818183C66666600;
            8'h5A : font_char = 64'h7F070E1C38707F00;
            8'h5B : font_char = 64'h3E06060606063E00;
            8'h5C : font_char = 64'h406030180C060200;
            8'h5D : font_char = 64'h3E30303030303E00;
            8'h5E : font_char = 64'h00000063361C0800;
            8'h5F : font_char = 64'h7F00000000000000;
            8'h60 : font_char = 64'h0000000000080400;
            8'h61 : font_char = 64'h7E637E603E000000;
            8'h62 : font_char = 64'h3F6363633F030300;
            8'h63 : font_char = 64'h3E6303633E000000;
            8'h64 : font_char = 64'h7E6363637E606000;
            8'h65 : font_char = 64'h3E037F633E000000;
            8'h66 : font_char = 64'h0C0C0C0C7F0C3C00;
            8'h67 : font_char = 64'h3E607E637E000000;
            8'h68 : font_char = 64'h636363633F030300;
            8'h69 : font_char = 64'h7F1818181E001800;
            8'h6A : font_char = 64'h3E63606060006000;
            8'h6B : font_char = 64'h63331F3363030300;
            8'h6C : font_char = 64'h780E030303030300;
            8'h6D : font_char = 64'h6B6B6B6B3F000000;
            8'h6E : font_char = 64'h636363633F000000;
            8'h6F : font_char = 64'h3E6363633E000000;
            8'h70 : font_char = 64'h03033F633F000000;
            8'h71 : font_char = 64'h60607E637E000000;
            8'h72 : font_char = 64'h030303673B000000;
            8'h73 : font_char = 64'h3F607F037E000000;
            8'h74 : font_char = 64'h7C0C0C0C7F0C0C00;
            8'h75 : font_char = 64'h3E63636363000000;
            8'h76 : font_char = 64'h081C366363000000;
            8'h77 : font_char = 64'h367F6B6B63000000;
            8'h78 : font_char = 64'h773E1C3E77000000;
            8'h79 : font_char = 64'h0F1C366363000000;
            8'h7A : font_char = 64'h7F0E1C387F000000;
            8'h7B : font_char = 64'h380C0C0E0C0C3800;
            8'h7C : font_char = 64'h0C0C0C0C0C0C0C00;
            8'h7D : font_char = 64'h0E18183818180E00;
            8'h7E : font_char = 64'h003B6B6E00000000;
            8'hA1 : font_char = 64'h0C1E1E1E0C000C00;
            8'hA2 : font_char = 64'h083E6B0B6B3E0800;
            8'hA3 : font_char = 64'h7F06061F46663C00;
            8'hA4 : font_char = 64'h00221C141C220000;
            8'hA5 : font_char = 64'h083E083E1C366300;
            8'hA6 : font_char = 64'h0C0C0C000C0C0C00;
            8'hA7 : font_char = 64'h3C607E633F031E00;
            8'hA8 : font_char = 64'h0000000000003600;
            8'hA9 : font_char = 64'h3E415D455D413E00;
            8'hAA : font_char = 64'h00007E637E603E00;
            8'hAB : font_char = 64'h6C361B366C000000;
            8'hAC : font_char = 64'h0030303E00000000;
            8'hAD : font_char = 64'h00003E0000000000;
            8'hAE : font_char = 64'h3E41454D55413E00;
            8'hAF : font_char = 64'h0000000000003E00;
            8'hB0 : font_char = 64'h00003E6763733E00;
            8'hB1 : font_char = 64'h3E0008083E080800;
            8'hB2 : font_char = 64'h00007E0C38633E00;
            8'hB3 : font_char = 64'h00003E6338633E00;
            8'hB4 : font_char = 64'h0000000000081000;
            8'hB5 : font_char = 64'h03033F6363636300;
            8'hB6 : font_char = 64'h28282C2E2F2E7C00;
            8'hB7 : font_char = 64'h0000000800000000;
            8'hB8 : font_char = 64'h0408000000000000;
            8'hB9 : font_char = 64'h00007E1818181E00;
            8'hBA : font_char = 64'h00003E6363633E00;
            8'hBB : font_char = 64'h1B366C361B000000;
            8'hBC : font_char = 64'h4040775252030200;
            8'hBD : font_char = 64'h7010274232030200;
            8'hBE : font_char = 64'h4040735452040300;
            8'hBF : font_char = 64'h3E63031E18001800;
            8'hC0 : font_char = 64'h637F63361C080400;
            8'hC1 : font_char = 64'h637F63361C081000;
            8'hC2 : font_char = 64'h637F63361C140800;
            8'hC3 : font_char = 64'h637F63361C142800;
            8'hC4 : font_char = 64'h637F63361C003600;
            8'hC5 : font_char = 64'h637F63361C141C00;
            8'hC6 : font_char = 64'h7B1B1F7B1B1E7C00;
            8'hC7 : font_char = 64'h04083E6303633E00;
            8'hC8 : font_char = 64'h7F031F037F080400;
            8'hC9 : font_char = 64'h7F031F037F081000;
            8'hCA : font_char = 64'h7F031F037F140800;
            8'hCB : font_char = 64'h7F031F037F003600;
            8'hCC : font_char = 64'h7F1C1C1C7F080400;
            8'hCD : font_char = 64'h7F1C1C1C7F081000;
            8'hCE : font_char = 64'h7F1C1C1C7F140800;
            8'hCF : font_char = 64'h7F1C1C1C7F003600;
            8'hD0 : font_char = 64'h1E36666F66361E00;
            8'hD1 : font_char = 64'h63736B6763142800;
            8'hD2 : font_char = 64'h3E6363633E080400;
            8'hD3 : font_char = 64'h3E6363633E081000;
            8'hD4 : font_char = 64'h3E6363633E140800;
            8'hD5 : font_char = 64'h3E6363633E142800;
            8'hD6 : font_char = 64'h3E6363633E003600;
            8'hD7 : font_char = 64'h2214081422000000;
            8'hD8 : font_char = 64'h3E63676B73633E00;
            8'hD9 : font_char = 64'h3E63636363080400;
            8'hDA : font_char = 64'h3E63636363081000;
            8'hDB : font_char = 64'h3E63636363140800;
            8'hDC : font_char = 64'h3E63636363003600;
            8'hDD : font_char = 64'h1C1C3E6363081000;
            8'hDE : font_char = 64'h033F6363633F0300;
            8'hDF : font_char = 64'h3B6B633B1B331E00;
            8'hE0 : font_char = 64'h7E637E603E080400;
            8'hE1 : font_char = 64'h7E637E603E081000;
            8'hE2 : font_char = 64'h7E637E603E140800;
            8'hE3 : font_char = 64'h7E637E603E142800;
            8'hE4 : font_char = 64'h7E637E603E003600;
            8'hE5 : font_char = 64'h7E637E603E141C00;
            8'hE6 : font_char = 64'h3F0D7F6C3F000000;
            8'hE7 : font_char = 64'h04087E03037E0000;
            8'hE8 : font_char = 64'h3E037F633E080400;
            8'hE9 : font_char = 64'h3E037F633E081000;
            8'hEA : font_char = 64'h3E037F633E140800;
            8'hEB : font_char = 64'h3E037F633E003600;
            8'hEC : font_char = 64'h7F1818181E080400;
            8'hED : font_char = 64'h7F1818181E081000;
            8'hEE : font_char = 64'h7F1818181E140800;
            8'hEF : font_char = 64'h7F1818181E003600;
            8'hF0 : font_char = 64'h3E6363637E301800;
            8'hF1 : font_char = 64'h636363633F142800;
            8'hF2 : font_char = 64'h3E63633E00080400;
            8'hF3 : font_char = 64'h3E63633E00081000;
            8'hF4 : font_char = 64'h3E63633E00140800;
            8'hF5 : font_char = 64'h3E63633E00142800;
            8'hF6 : font_char = 64'h3E63633E00360000;
            8'hF7 : font_char = 64'h08003E0008000000;
            8'hF8 : font_char = 64'h3E676B733E000000;
            8'hF9 : font_char = 64'h3E63636300080400;
            8'hFA : font_char = 64'h3E63636300081000;
            8'hFB : font_char = 64'h3E63636300140800;
            8'hFC : font_char = 64'h3E63636300360000;
            8'hFD : font_char = 64'h0F1C366363081000;
            8'hFE : font_char = 64'h03033F633F030300;
            8'hFF : font_char = 64'h0F1C366363003600;
            default : font_char = 64'h0;
        endcase

endmodule

