
module reflet_VGA_txt #(
    parameter h_size = 640,
    v_size = 480,
    color_depth = 8,


